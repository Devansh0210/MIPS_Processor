module RegFile(
      input wire[3:0] inp_add,
      output wire out_add
);



endmodule